	component lab is
	end component lab;

	u0 : component lab
		port map (
		);

