-- lab1_system.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lab1_system is
	port (
		hps_io_hps_io_usb1_inst_D0  : inout std_logic                     := '0';             --               hps_io.hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1  : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2  : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3  : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4  : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5  : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6  : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7  : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK : in    std_logic                     := '0';             --                     .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP : out   std_logic;                                        --                     .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR : in    std_logic                     := '0';             --                     .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT : in    std_logic                     := '0';             --                     .hps_io_usb1_inst_NXT
		hps_io_hps_io_uart0_inst_RX : in    std_logic                     := '0';             --                     .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX : out   std_logic;                                        --                     .hps_io_uart0_inst_TX
		leds_readdata               : out   std_logic_vector(9 downto 0);                     --                 leds.readdata
		memory_mem_a                : out   std_logic_vector(14 downto 0);                    --               memory.mem_a
		memory_mem_ba               : out   std_logic_vector(2 downto 0);                     --                     .mem_ba
		memory_mem_ck               : out   std_logic;                                        --                     .mem_ck
		memory_mem_ck_n             : out   std_logic;                                        --                     .mem_ck_n
		memory_mem_cke              : out   std_logic;                                        --                     .mem_cke
		memory_mem_cs_n             : out   std_logic;                                        --                     .mem_cs_n
		memory_mem_ras_n            : out   std_logic;                                        --                     .mem_ras_n
		memory_mem_cas_n            : out   std_logic;                                        --                     .mem_cas_n
		memory_mem_we_n             : out   std_logic;                                        --                     .mem_we_n
		memory_mem_reset_n          : out   std_logic;                                        --                     .mem_reset_n
		memory_mem_dq               : inout std_logic_vector(31 downto 0) := (others => '0'); --                     .mem_dq
		memory_mem_dqs              : inout std_logic_vector(3 downto 0)  := (others => '0'); --                     .mem_dqs
		memory_mem_dqs_n            : inout std_logic_vector(3 downto 0)  := (others => '0'); --                     .mem_dqs_n
		memory_mem_odt              : out   std_logic;                                        --                     .mem_odt
		memory_mem_dm               : out   std_logic_vector(3 downto 0);                     --                     .mem_dm
		memory_oct_rzqin            : in    std_logic                     := '0';             --                     .oct_rzqin
		pushbuttons_export          : in    std_logic_vector(3 downto 0)  := (others => '0'); --          pushbuttons.export
		system_pll_ref_clk_clk      : in    std_logic                     := '0';             --   system_pll_ref_clk.clk
		system_pll_ref_reset_reset  : in    std_logic                     := '0'              -- system_pll_ref_reset.reset
	);
end entity lab1_system;

architecture rtl of lab1_system is
	component lab1_system_ARM_A9_HPS is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			f2h_stm_hwevents     : in    std_logic_vector(27 downto 0) := (others => 'X'); -- stm_hwevents
			mem_a                : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba               : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck               : out   std_logic;                                        -- mem_ck
			mem_ck_n             : out   std_logic;                                        -- mem_ck_n
			mem_cke              : out   std_logic;                                        -- mem_cke
			mem_cs_n             : out   std_logic;                                        -- mem_cs_n
			mem_ras_n            : out   std_logic;                                        -- mem_ras_n
			mem_cas_n            : out   std_logic;                                        -- mem_cas_n
			mem_we_n             : out   std_logic;                                        -- mem_we_n
			mem_reset_n          : out   std_logic;                                        -- mem_reset_n
			mem_dq               : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs              : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n            : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt              : out   std_logic;                                        -- mem_odt
			mem_dm               : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin            : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_usb1_inst_D0  : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1  : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2  : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3  : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4  : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5  : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6  : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7  : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_uart0_inst_RX : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX : out   std_logic;                                        -- hps_io_uart0_inst_TX
			h2f_rst_n            : out   std_logic;                                        -- reset_n
			h2f_axi_clk          : in    std_logic                     := 'X';             -- clk
			h2f_AWID             : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR           : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN            : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE           : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST          : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK           : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE          : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT           : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID          : out   std_logic;                                        -- awvalid
			h2f_AWREADY          : in    std_logic                     := 'X';             -- awready
			h2f_WID              : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA            : out   std_logic_vector(63 downto 0);                    -- wdata
			h2f_WSTRB            : out   std_logic_vector(7 downto 0);                     -- wstrb
			h2f_WLAST            : out   std_logic;                                        -- wlast
			h2f_WVALID           : out   std_logic;                                        -- wvalid
			h2f_WREADY           : in    std_logic                     := 'X';             -- wready
			h2f_BID              : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP            : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID           : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY           : out   std_logic;                                        -- bready
			h2f_ARID             : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR           : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN            : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE           : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST          : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK           : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE          : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT           : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID          : out   std_logic;                                        -- arvalid
			h2f_ARREADY          : in    std_logic                     := 'X';             -- arready
			h2f_RID              : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA            : in    std_logic_vector(63 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP            : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST            : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID           : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY           : out   std_logic;                                        -- rready
			f2h_axi_clk          : in    std_logic                     := 'X';             -- clk
			f2h_AWID             : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- awid
			f2h_AWADDR           : in    std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			f2h_AWLEN            : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			f2h_AWSIZE           : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			f2h_AWBURST          : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			f2h_AWLOCK           : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			f2h_AWCACHE          : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			f2h_AWPROT           : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			f2h_AWVALID          : in    std_logic                     := 'X';             -- awvalid
			f2h_AWREADY          : out   std_logic;                                        -- awready
			f2h_AWUSER           : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- awuser
			f2h_WID              : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wid
			f2h_WDATA            : in    std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB            : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST            : in    std_logic                     := 'X';             -- wlast
			f2h_WVALID           : in    std_logic                     := 'X';             -- wvalid
			f2h_WREADY           : out   std_logic;                                        -- wready
			f2h_BID              : out   std_logic_vector(7 downto 0);                     -- bid
			f2h_BRESP            : out   std_logic_vector(1 downto 0);                     -- bresp
			f2h_BVALID           : out   std_logic;                                        -- bvalid
			f2h_BREADY           : in    std_logic                     := 'X';             -- bready
			f2h_ARID             : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- arid
			f2h_ARADDR           : in    std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			f2h_ARLEN            : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			f2h_ARSIZE           : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			f2h_ARBURST          : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			f2h_ARLOCK           : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			f2h_ARCACHE          : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			f2h_ARPROT           : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			f2h_ARVALID          : in    std_logic                     := 'X';             -- arvalid
			f2h_ARREADY          : out   std_logic;                                        -- arready
			f2h_ARUSER           : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- aruser
			f2h_RID              : out   std_logic_vector(7 downto 0);                     -- rid
			f2h_RDATA            : out   std_logic_vector(63 downto 0);                    -- rdata
			f2h_RRESP            : out   std_logic_vector(1 downto 0);                     -- rresp
			f2h_RLAST            : out   std_logic;                                        -- rlast
			f2h_RVALID           : out   std_logic;                                        -- rvalid
			f2h_RREADY           : in    std_logic                     := 'X';             -- rready
			h2f_lw_axi_clk       : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID          : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR        : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN         : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE        : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST       : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK        : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE       : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT        : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID       : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY       : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID           : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA         : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB         : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST         : out   std_logic;                                        -- wlast
			h2f_lw_WVALID        : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY        : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID           : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP         : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID        : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY        : out   std_logic;                                        -- bready
			h2f_lw_ARID          : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR        : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN         : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE        : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST       : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK        : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE       : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT        : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID       : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY       : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID           : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA         : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP         : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST         : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID        : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY        : out   std_logic;                                        -- rready
			f2h_irq_p0           : in    std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			f2h_irq_p1           : in    std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component lab1_system_ARM_A9_HPS;

	component lab1_system_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component lab1_system_JTAG_UART;

	component lab1_system_Pushbuttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component lab1_system_Pushbuttons;

	component lab1_system_System_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component lab1_system_System_PLL;

	component axi4_lite_count28 is
		generic (
			C_S_AXI_DATA_WIDTH : integer := 32;
			C_S_AXI_ADDR_WIDTH : integer := 4
		);
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset_n            : in  std_logic                     := 'X';             -- reset_n
			out_leds           : out std_logic_vector(9 downto 0);                     -- readdata
			axs_s0_AXI_AWADDR  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awaddr
			axs_s0_AXI_AWPROT  : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			axs_s0_AXI_AWVALID : in  std_logic                     := 'X';             -- awvalid
			axs_s0_AXI_AWREADY : out std_logic;                                        -- awready
			axs_s0_AXI_WDATA   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			axs_s0_AXI_WSTRB   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			axs_s0_AXI_WVALID  : in  std_logic                     := 'X';             -- wvalid
			axs_s0_AXI_WREADY  : out std_logic;                                        -- wready
			axs_s0_AXI_BRESP   : out std_logic_vector(1 downto 0);                     -- bresp
			axs_s0_AXI_BVALID  : out std_logic;                                        -- bvalid
			axs_s0_AXI_BREADY  : in  std_logic                     := 'X';             -- bready
			axs_s0_AXI_ARADDR  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- araddr
			axs_s0_AXI_ARPROT  : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			axs_s0_AXI_ARVALID : in  std_logic                     := 'X';             -- arvalid
			axs_s0_AXI_ARREADY : out std_logic;                                        -- arready
			axs_s0_AXI_RDATA   : out std_logic_vector(31 downto 0);                    -- rdata
			axs_s0_AXI_RRESP   : out std_logic_vector(1 downto 0);                     -- rresp
			axs_s0_AXI_RVALID  : out std_logic;                                        -- rvalid
			axs_s0_AXI_RREADY  : in  std_logic                     := 'X'              -- rready
		);
	end component axi4_lite_count28;

	component lab1_system_mm_interconnect_0 is
		port (
			ARM_A9_HPS_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			ARM_A9_HPS_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			ARM_A9_HPS_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			ARM_A9_HPS_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			ARM_A9_HPS_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			ARM_A9_HPS_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			ARM_A9_HPS_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			ARM_A9_HPS_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			ARM_A9_HPS_h2f_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			ARM_A9_HPS_h2f_axi_master_awready                                     : out std_logic;                                        -- awready
			ARM_A9_HPS_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			ARM_A9_HPS_h2f_axi_master_wdata                                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			ARM_A9_HPS_h2f_axi_master_wstrb                                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			ARM_A9_HPS_h2f_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			ARM_A9_HPS_h2f_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			ARM_A9_HPS_h2f_axi_master_wready                                      : out std_logic;                                        -- wready
			ARM_A9_HPS_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			ARM_A9_HPS_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			ARM_A9_HPS_h2f_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			ARM_A9_HPS_h2f_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			ARM_A9_HPS_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			ARM_A9_HPS_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			ARM_A9_HPS_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			ARM_A9_HPS_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			ARM_A9_HPS_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			ARM_A9_HPS_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			ARM_A9_HPS_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			ARM_A9_HPS_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			ARM_A9_HPS_h2f_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			ARM_A9_HPS_h2f_axi_master_arready                                     : out std_logic;                                        -- arready
			ARM_A9_HPS_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			ARM_A9_HPS_h2f_axi_master_rdata                                       : out std_logic_vector(63 downto 0);                    -- rdata
			ARM_A9_HPS_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			ARM_A9_HPS_h2f_axi_master_rlast                                       : out std_logic;                                        -- rlast
			ARM_A9_HPS_h2f_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			ARM_A9_HPS_h2f_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			System_PLL_sys_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			JTAG_UART_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			JTAG_UART_avalon_jtag_slave_address                                   : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write                                     : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read                                      : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect                                : out std_logic                                         -- chipselect
		);
	end component lab1_system_mm_interconnect_0;

	component lab1_system_mm_interconnect_1 is
		port (
			ARM_A9_HPS_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			ARM_A9_HPS_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			ARM_A9_HPS_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			ARM_A9_HPS_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			ARM_A9_HPS_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			ARM_A9_HPS_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			ARM_A9_HPS_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			ARM_A9_HPS_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			ARM_A9_HPS_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			ARM_A9_HPS_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			ARM_A9_HPS_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			ARM_A9_HPS_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			ARM_A9_HPS_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			ARM_A9_HPS_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			ARM_A9_HPS_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			ARM_A9_HPS_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			ARM_A9_HPS_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			ARM_A9_HPS_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			ARM_A9_HPS_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			ARM_A9_HPS_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			ARM_A9_HPS_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			ARM_A9_HPS_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			ARM_A9_HPS_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			ARM_A9_HPS_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			ARM_A9_HPS_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			ARM_A9_HPS_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			ARM_A9_HPS_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			ARM_A9_HPS_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			ARM_A9_HPS_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			axi4_lite_count28_0_axi4_lite_awaddr                                     : out std_logic_vector(3 downto 0);                     -- awaddr
			axi4_lite_count28_0_axi4_lite_awprot                                     : out std_logic_vector(2 downto 0);                     -- awprot
			axi4_lite_count28_0_axi4_lite_awvalid                                    : out std_logic;                                        -- awvalid
			axi4_lite_count28_0_axi4_lite_awready                                    : in  std_logic                     := 'X';             -- awready
			axi4_lite_count28_0_axi4_lite_wdata                                      : out std_logic_vector(31 downto 0);                    -- wdata
			axi4_lite_count28_0_axi4_lite_wstrb                                      : out std_logic_vector(3 downto 0);                     -- wstrb
			axi4_lite_count28_0_axi4_lite_wvalid                                     : out std_logic;                                        -- wvalid
			axi4_lite_count28_0_axi4_lite_wready                                     : in  std_logic                     := 'X';             -- wready
			axi4_lite_count28_0_axi4_lite_bresp                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			axi4_lite_count28_0_axi4_lite_bvalid                                     : in  std_logic                     := 'X';             -- bvalid
			axi4_lite_count28_0_axi4_lite_bready                                     : out std_logic;                                        -- bready
			axi4_lite_count28_0_axi4_lite_araddr                                     : out std_logic_vector(3 downto 0);                     -- araddr
			axi4_lite_count28_0_axi4_lite_arprot                                     : out std_logic_vector(2 downto 0);                     -- arprot
			axi4_lite_count28_0_axi4_lite_arvalid                                    : out std_logic;                                        -- arvalid
			axi4_lite_count28_0_axi4_lite_arready                                    : in  std_logic                     := 'X';             -- arready
			axi4_lite_count28_0_axi4_lite_rdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			axi4_lite_count28_0_axi4_lite_rresp                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			axi4_lite_count28_0_axi4_lite_rvalid                                     : in  std_logic                     := 'X';             -- rvalid
			axi4_lite_count28_0_axi4_lite_rready                                     : out std_logic;                                        -- rready
			System_PLL_sys_clk_clk                                                   : in  std_logic                     := 'X';             -- clk
			ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			axi4_lite_count28_0_reset_reset_bridge_in_reset_reset                    : in  std_logic                     := 'X';             -- reset
			Pushbuttons_reset_reset_bridge_in_reset_reset                            : in  std_logic                     := 'X';             -- reset
			Pushbuttons_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			Pushbuttons_s1_write                                                     : out std_logic;                                        -- write
			Pushbuttons_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Pushbuttons_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			Pushbuttons_s1_chipselect                                                : out std_logic                                         -- chipselect
		);
	end component lab1_system_mm_interconnect_1;

	component lab1_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component lab1_system_irq_mapper;

	component lab1_system_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component lab1_system_irq_mapper_001;

	component lab1_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab1_system_rst_controller;

	component lab1_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab1_system_rst_controller_001;

	signal system_pll_sys_clk_clk                                        : std_logic;                     -- System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, JTAG_UART:clk, Pushbuttons:clk, axi4_lite_count28_0:clk, mm_interconnect_0:System_PLL_sys_clk_clk, mm_interconnect_1:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk]
	signal arm_a9_hps_h2f_axi_master_awburst                             : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awburst
	signal arm_a9_hps_h2f_axi_master_arlen                               : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlen
	signal arm_a9_hps_h2f_axi_master_wstrb                               : std_logic_vector(7 downto 0);  -- ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wstrb
	signal arm_a9_hps_h2f_axi_master_wready                              : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	signal arm_a9_hps_h2f_axi_master_rid                                 : std_logic_vector(11 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	signal arm_a9_hps_h2f_axi_master_rready                              : std_logic;                     -- ARM_A9_HPS:h2f_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rready
	signal arm_a9_hps_h2f_axi_master_awlen                               : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlen
	signal arm_a9_hps_h2f_axi_master_wid                                 : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wid
	signal arm_a9_hps_h2f_axi_master_arcache                             : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arcache
	signal arm_a9_hps_h2f_axi_master_wvalid                              : std_logic;                     -- ARM_A9_HPS:h2f_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wvalid
	signal arm_a9_hps_h2f_axi_master_araddr                              : std_logic_vector(29 downto 0); -- ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_araddr
	signal arm_a9_hps_h2f_axi_master_arprot                              : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arprot
	signal arm_a9_hps_h2f_axi_master_awprot                              : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awprot
	signal arm_a9_hps_h2f_axi_master_wdata                               : std_logic_vector(63 downto 0); -- ARM_A9_HPS:h2f_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wdata
	signal arm_a9_hps_h2f_axi_master_arvalid                             : std_logic;                     -- ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arvalid
	signal arm_a9_hps_h2f_axi_master_awcache                             : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awcache
	signal arm_a9_hps_h2f_axi_master_arid                                : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arid
	signal arm_a9_hps_h2f_axi_master_arlock                              : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlock
	signal arm_a9_hps_h2f_axi_master_awlock                              : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlock
	signal arm_a9_hps_h2f_axi_master_awaddr                              : std_logic_vector(29 downto 0); -- ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awaddr
	signal arm_a9_hps_h2f_axi_master_bresp                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	signal arm_a9_hps_h2f_axi_master_arready                             : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	signal arm_a9_hps_h2f_axi_master_rdata                               : std_logic_vector(63 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	signal arm_a9_hps_h2f_axi_master_awready                             : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	signal arm_a9_hps_h2f_axi_master_arburst                             : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arburst
	signal arm_a9_hps_h2f_axi_master_arsize                              : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arsize
	signal arm_a9_hps_h2f_axi_master_bready                              : std_logic;                     -- ARM_A9_HPS:h2f_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bready
	signal arm_a9_hps_h2f_axi_master_rlast                               : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	signal arm_a9_hps_h2f_axi_master_wlast                               : std_logic;                     -- ARM_A9_HPS:h2f_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wlast
	signal arm_a9_hps_h2f_axi_master_rresp                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	signal arm_a9_hps_h2f_axi_master_awid                                : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awid
	signal arm_a9_hps_h2f_axi_master_bid                                 : std_logic_vector(11 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	signal arm_a9_hps_h2f_axi_master_bvalid                              : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	signal arm_a9_hps_h2f_axi_master_awsize                              : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awsize
	signal arm_a9_hps_h2f_axi_master_awvalid                             : std_logic;                     -- ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awvalid
	signal arm_a9_hps_h2f_axi_master_rvalid                              : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal arm_a9_hps_h2f_lw_axi_master_awburst                          : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awburst
	signal arm_a9_hps_h2f_lw_axi_master_arlen                            : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arlen
	signal arm_a9_hps_h2f_lw_axi_master_wstrb                            : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	signal arm_a9_hps_h2f_lw_axi_master_wready                           : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	signal arm_a9_hps_h2f_lw_axi_master_rid                              : std_logic_vector(11 downto 0); -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	signal arm_a9_hps_h2f_lw_axi_master_rready                           : std_logic;                     -- ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rready
	signal arm_a9_hps_h2f_lw_axi_master_awlen                            : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awlen
	signal arm_a9_hps_h2f_lw_axi_master_wid                              : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wid
	signal arm_a9_hps_h2f_lw_axi_master_arcache                          : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arcache
	signal arm_a9_hps_h2f_lw_axi_master_wvalid                           : std_logic;                     -- ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	signal arm_a9_hps_h2f_lw_axi_master_araddr                           : std_logic_vector(20 downto 0); -- ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_araddr
	signal arm_a9_hps_h2f_lw_axi_master_arprot                           : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arprot
	signal arm_a9_hps_h2f_lw_axi_master_awprot                           : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awprot
	signal arm_a9_hps_h2f_lw_axi_master_wdata                            : std_logic_vector(31 downto 0); -- ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wdata
	signal arm_a9_hps_h2f_lw_axi_master_arvalid                          : std_logic;                     -- ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	signal arm_a9_hps_h2f_lw_axi_master_awcache                          : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awcache
	signal arm_a9_hps_h2f_lw_axi_master_arid                             : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arid
	signal arm_a9_hps_h2f_lw_axi_master_arlock                           : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arlock
	signal arm_a9_hps_h2f_lw_axi_master_awlock                           : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awlock
	signal arm_a9_hps_h2f_lw_axi_master_awaddr                           : std_logic_vector(20 downto 0); -- ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	signal arm_a9_hps_h2f_lw_axi_master_bresp                            : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	signal arm_a9_hps_h2f_lw_axi_master_arready                          : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	signal arm_a9_hps_h2f_lw_axi_master_rdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	signal arm_a9_hps_h2f_lw_axi_master_awready                          : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	signal arm_a9_hps_h2f_lw_axi_master_arburst                          : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arburst
	signal arm_a9_hps_h2f_lw_axi_master_arsize                           : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arsize
	signal arm_a9_hps_h2f_lw_axi_master_bready                           : std_logic;                     -- ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bready
	signal arm_a9_hps_h2f_lw_axi_master_rlast                            : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	signal arm_a9_hps_h2f_lw_axi_master_wlast                            : std_logic;                     -- ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wlast
	signal arm_a9_hps_h2f_lw_axi_master_rresp                            : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	signal arm_a9_hps_h2f_lw_axi_master_awid                             : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awid
	signal arm_a9_hps_h2f_lw_axi_master_bid                              : std_logic_vector(11 downto 0); -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	signal arm_a9_hps_h2f_lw_axi_master_bvalid                           : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	signal arm_a9_hps_h2f_lw_axi_master_awsize                           : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awsize
	signal arm_a9_hps_h2f_lw_axi_master_awvalid                          : std_logic;                     -- ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	signal arm_a9_hps_h2f_lw_axi_master_rvalid                           : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awaddr        : std_logic_vector(3 downto 0);  -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_awaddr -> axi4_lite_count28_0:axs_s0_AXI_AWADDR
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bresp         : std_logic_vector(1 downto 0);  -- axi4_lite_count28_0:axs_s0_AXI_BRESP -> mm_interconnect_1:axi4_lite_count28_0_axi4_lite_bresp
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arready       : std_logic;                     -- axi4_lite_count28_0:axs_s0_AXI_ARREADY -> mm_interconnect_1:axi4_lite_count28_0_axi4_lite_arready
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rdata         : std_logic_vector(31 downto 0); -- axi4_lite_count28_0:axs_s0_AXI_RDATA -> mm_interconnect_1:axi4_lite_count28_0_axi4_lite_rdata
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wstrb         : std_logic_vector(3 downto 0);  -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_wstrb -> axi4_lite_count28_0:axs_s0_AXI_WSTRB
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wready        : std_logic;                     -- axi4_lite_count28_0:axs_s0_AXI_WREADY -> mm_interconnect_1:axi4_lite_count28_0_axi4_lite_wready
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awready       : std_logic;                     -- axi4_lite_count28_0:axs_s0_AXI_AWREADY -> mm_interconnect_1:axi4_lite_count28_0_axi4_lite_awready
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rready        : std_logic;                     -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_rready -> axi4_lite_count28_0:axs_s0_AXI_RREADY
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bready        : std_logic;                     -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_bready -> axi4_lite_count28_0:axs_s0_AXI_BREADY
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wvalid        : std_logic;                     -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_wvalid -> axi4_lite_count28_0:axs_s0_AXI_WVALID
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_araddr        : std_logic_vector(3 downto 0);  -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_araddr -> axi4_lite_count28_0:axs_s0_AXI_ARADDR
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arprot        : std_logic_vector(2 downto 0);  -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_arprot -> axi4_lite_count28_0:axs_s0_AXI_ARPROT
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rresp         : std_logic_vector(1 downto 0);  -- axi4_lite_count28_0:axs_s0_AXI_RRESP -> mm_interconnect_1:axi4_lite_count28_0_axi4_lite_rresp
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awprot        : std_logic_vector(2 downto 0);  -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_awprot -> axi4_lite_count28_0:axs_s0_AXI_AWPROT
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wdata         : std_logic_vector(31 downto 0); -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_wdata -> axi4_lite_count28_0:axs_s0_AXI_WDATA
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arvalid       : std_logic;                     -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_arvalid -> axi4_lite_count28_0:axs_s0_AXI_ARVALID
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bvalid        : std_logic;                     -- axi4_lite_count28_0:axs_s0_AXI_BVALID -> mm_interconnect_1:axi4_lite_count28_0_axi4_lite_bvalid
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awvalid       : std_logic;                     -- mm_interconnect_1:axi4_lite_count28_0_axi4_lite_awvalid -> axi4_lite_count28_0:axs_s0_AXI_AWVALID
	signal mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rvalid        : std_logic;                     -- axi4_lite_count28_0:axs_s0_AXI_RVALID -> mm_interconnect_1:axi4_lite_count28_0_axi4_lite_rvalid
	signal mm_interconnect_1_pushbuttons_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:Pushbuttons_s1_chipselect -> Pushbuttons:chipselect
	signal mm_interconnect_1_pushbuttons_s1_readdata                     : std_logic_vector(31 downto 0); -- Pushbuttons:readdata -> mm_interconnect_1:Pushbuttons_s1_readdata
	signal mm_interconnect_1_pushbuttons_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:Pushbuttons_s1_address -> Pushbuttons:address
	signal mm_interconnect_1_pushbuttons_s1_write                        : std_logic;                     -- mm_interconnect_1:Pushbuttons_s1_write -> mm_interconnect_1_pushbuttons_s1_write:in
	signal mm_interconnect_1_pushbuttons_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:Pushbuttons_s1_writedata -> Pushbuttons:writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- Pushbuttons:irq -> irq_mapper:receiver1_irq
	signal arm_a9_hps_f2h_irq0_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	signal arm_a9_hps_f2h_irq1_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:JTAG_UART_reset_reset_bridge_in_reset_reset, mm_interconnect_1:axi4_lite_count28_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal arm_a9_hps_h2f_reset_reset                                    : std_logic;                     -- ARM_A9_HPS:h2f_rst_n -> arm_a9_hps_h2f_reset_reset:in
	signal system_pll_reset_source_reset                                 : std_logic;                     -- System_PLL:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_1:Pushbuttons_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_1_pushbuttons_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_1_pushbuttons_s1_write:inv -> Pushbuttons:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [JTAG_UART:rst_n, axi4_lite_count28_0:reset_n]
	signal arm_a9_hps_h2f_reset_reset_ports_inv                          : std_logic;                     -- arm_a9_hps_h2f_reset_reset:inv -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> Pushbuttons:reset_n

begin

	arm_a9_hps : component lab1_system_ARM_A9_HPS
		generic map (
			F2S_Width => 2,
			S2F_Width => 2
		)
		port map (
			f2h_stm_hwevents     => open,                                 -- f2h_stm_hw_events.stm_hwevents
			mem_a                => memory_mem_a,                         --            memory.mem_a
			mem_ba               => memory_mem_ba,                        --                  .mem_ba
			mem_ck               => memory_mem_ck,                        --                  .mem_ck
			mem_ck_n             => memory_mem_ck_n,                      --                  .mem_ck_n
			mem_cke              => memory_mem_cke,                       --                  .mem_cke
			mem_cs_n             => memory_mem_cs_n,                      --                  .mem_cs_n
			mem_ras_n            => memory_mem_ras_n,                     --                  .mem_ras_n
			mem_cas_n            => memory_mem_cas_n,                     --                  .mem_cas_n
			mem_we_n             => memory_mem_we_n,                      --                  .mem_we_n
			mem_reset_n          => memory_mem_reset_n,                   --                  .mem_reset_n
			mem_dq               => memory_mem_dq,                        --                  .mem_dq
			mem_dqs              => memory_mem_dqs,                       --                  .mem_dqs
			mem_dqs_n            => memory_mem_dqs_n,                     --                  .mem_dqs_n
			mem_odt              => memory_mem_odt,                       --                  .mem_odt
			mem_dm               => memory_mem_dm,                        --                  .mem_dm
			oct_rzqin            => memory_oct_rzqin,                     --                  .oct_rzqin
			hps_io_usb1_inst_D0  => hps_io_hps_io_usb1_inst_D0,           --            hps_io.hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1  => hps_io_hps_io_usb1_inst_D1,           --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2  => hps_io_hps_io_usb1_inst_D2,           --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3  => hps_io_hps_io_usb1_inst_D3,           --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4  => hps_io_hps_io_usb1_inst_D4,           --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5  => hps_io_hps_io_usb1_inst_D5,           --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6  => hps_io_hps_io_usb1_inst_D6,           --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7  => hps_io_hps_io_usb1_inst_D7,           --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK => hps_io_hps_io_usb1_inst_CLK,          --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP => hps_io_hps_io_usb1_inst_STP,          --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR => hps_io_hps_io_usb1_inst_DIR,          --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT => hps_io_hps_io_usb1_inst_NXT,          --                  .hps_io_usb1_inst_NXT
			hps_io_uart0_inst_RX => hps_io_hps_io_uart0_inst_RX,          --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX => hps_io_hps_io_uart0_inst_TX,          --                  .hps_io_uart0_inst_TX
			h2f_rst_n            => arm_a9_hps_h2f_reset_reset,           --         h2f_reset.reset_n
			h2f_axi_clk          => system_pll_sys_clk_clk,               --     h2f_axi_clock.clk
			h2f_AWID             => arm_a9_hps_h2f_axi_master_awid,       --    h2f_axi_master.awid
			h2f_AWADDR           => arm_a9_hps_h2f_axi_master_awaddr,     --                  .awaddr
			h2f_AWLEN            => arm_a9_hps_h2f_axi_master_awlen,      --                  .awlen
			h2f_AWSIZE           => arm_a9_hps_h2f_axi_master_awsize,     --                  .awsize
			h2f_AWBURST          => arm_a9_hps_h2f_axi_master_awburst,    --                  .awburst
			h2f_AWLOCK           => arm_a9_hps_h2f_axi_master_awlock,     --                  .awlock
			h2f_AWCACHE          => arm_a9_hps_h2f_axi_master_awcache,    --                  .awcache
			h2f_AWPROT           => arm_a9_hps_h2f_axi_master_awprot,     --                  .awprot
			h2f_AWVALID          => arm_a9_hps_h2f_axi_master_awvalid,    --                  .awvalid
			h2f_AWREADY          => arm_a9_hps_h2f_axi_master_awready,    --                  .awready
			h2f_WID              => arm_a9_hps_h2f_axi_master_wid,        --                  .wid
			h2f_WDATA            => arm_a9_hps_h2f_axi_master_wdata,      --                  .wdata
			h2f_WSTRB            => arm_a9_hps_h2f_axi_master_wstrb,      --                  .wstrb
			h2f_WLAST            => arm_a9_hps_h2f_axi_master_wlast,      --                  .wlast
			h2f_WVALID           => arm_a9_hps_h2f_axi_master_wvalid,     --                  .wvalid
			h2f_WREADY           => arm_a9_hps_h2f_axi_master_wready,     --                  .wready
			h2f_BID              => arm_a9_hps_h2f_axi_master_bid,        --                  .bid
			h2f_BRESP            => arm_a9_hps_h2f_axi_master_bresp,      --                  .bresp
			h2f_BVALID           => arm_a9_hps_h2f_axi_master_bvalid,     --                  .bvalid
			h2f_BREADY           => arm_a9_hps_h2f_axi_master_bready,     --                  .bready
			h2f_ARID             => arm_a9_hps_h2f_axi_master_arid,       --                  .arid
			h2f_ARADDR           => arm_a9_hps_h2f_axi_master_araddr,     --                  .araddr
			h2f_ARLEN            => arm_a9_hps_h2f_axi_master_arlen,      --                  .arlen
			h2f_ARSIZE           => arm_a9_hps_h2f_axi_master_arsize,     --                  .arsize
			h2f_ARBURST          => arm_a9_hps_h2f_axi_master_arburst,    --                  .arburst
			h2f_ARLOCK           => arm_a9_hps_h2f_axi_master_arlock,     --                  .arlock
			h2f_ARCACHE          => arm_a9_hps_h2f_axi_master_arcache,    --                  .arcache
			h2f_ARPROT           => arm_a9_hps_h2f_axi_master_arprot,     --                  .arprot
			h2f_ARVALID          => arm_a9_hps_h2f_axi_master_arvalid,    --                  .arvalid
			h2f_ARREADY          => arm_a9_hps_h2f_axi_master_arready,    --                  .arready
			h2f_RID              => arm_a9_hps_h2f_axi_master_rid,        --                  .rid
			h2f_RDATA            => arm_a9_hps_h2f_axi_master_rdata,      --                  .rdata
			h2f_RRESP            => arm_a9_hps_h2f_axi_master_rresp,      --                  .rresp
			h2f_RLAST            => arm_a9_hps_h2f_axi_master_rlast,      --                  .rlast
			h2f_RVALID           => arm_a9_hps_h2f_axi_master_rvalid,     --                  .rvalid
			h2f_RREADY           => arm_a9_hps_h2f_axi_master_rready,     --                  .rready
			f2h_axi_clk          => system_pll_sys_clk_clk,               --     f2h_axi_clock.clk
			f2h_AWID             => open,                                 --     f2h_axi_slave.awid
			f2h_AWADDR           => open,                                 --                  .awaddr
			f2h_AWLEN            => open,                                 --                  .awlen
			f2h_AWSIZE           => open,                                 --                  .awsize
			f2h_AWBURST          => open,                                 --                  .awburst
			f2h_AWLOCK           => open,                                 --                  .awlock
			f2h_AWCACHE          => open,                                 --                  .awcache
			f2h_AWPROT           => open,                                 --                  .awprot
			f2h_AWVALID          => open,                                 --                  .awvalid
			f2h_AWREADY          => open,                                 --                  .awready
			f2h_AWUSER           => open,                                 --                  .awuser
			f2h_WID              => open,                                 --                  .wid
			f2h_WDATA            => open,                                 --                  .wdata
			f2h_WSTRB            => open,                                 --                  .wstrb
			f2h_WLAST            => open,                                 --                  .wlast
			f2h_WVALID           => open,                                 --                  .wvalid
			f2h_WREADY           => open,                                 --                  .wready
			f2h_BID              => open,                                 --                  .bid
			f2h_BRESP            => open,                                 --                  .bresp
			f2h_BVALID           => open,                                 --                  .bvalid
			f2h_BREADY           => open,                                 --                  .bready
			f2h_ARID             => open,                                 --                  .arid
			f2h_ARADDR           => open,                                 --                  .araddr
			f2h_ARLEN            => open,                                 --                  .arlen
			f2h_ARSIZE           => open,                                 --                  .arsize
			f2h_ARBURST          => open,                                 --                  .arburst
			f2h_ARLOCK           => open,                                 --                  .arlock
			f2h_ARCACHE          => open,                                 --                  .arcache
			f2h_ARPROT           => open,                                 --                  .arprot
			f2h_ARVALID          => open,                                 --                  .arvalid
			f2h_ARREADY          => open,                                 --                  .arready
			f2h_ARUSER           => open,                                 --                  .aruser
			f2h_RID              => open,                                 --                  .rid
			f2h_RDATA            => open,                                 --                  .rdata
			f2h_RRESP            => open,                                 --                  .rresp
			f2h_RLAST            => open,                                 --                  .rlast
			f2h_RVALID           => open,                                 --                  .rvalid
			f2h_RREADY           => open,                                 --                  .rready
			h2f_lw_axi_clk       => system_pll_sys_clk_clk,               --  h2f_lw_axi_clock.clk
			h2f_lw_AWID          => arm_a9_hps_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR        => arm_a9_hps_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN         => arm_a9_hps_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE        => arm_a9_hps_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST       => arm_a9_hps_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK        => arm_a9_hps_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE       => arm_a9_hps_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT        => arm_a9_hps_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID       => arm_a9_hps_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY       => arm_a9_hps_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID           => arm_a9_hps_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA         => arm_a9_hps_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB         => arm_a9_hps_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST         => arm_a9_hps_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID        => arm_a9_hps_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY        => arm_a9_hps_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID           => arm_a9_hps_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP         => arm_a9_hps_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID        => arm_a9_hps_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY        => arm_a9_hps_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID          => arm_a9_hps_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR        => arm_a9_hps_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN         => arm_a9_hps_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE        => arm_a9_hps_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST       => arm_a9_hps_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK        => arm_a9_hps_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE       => arm_a9_hps_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT        => arm_a9_hps_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID       => arm_a9_hps_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY       => arm_a9_hps_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID           => arm_a9_hps_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA         => arm_a9_hps_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP         => arm_a9_hps_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST         => arm_a9_hps_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID        => arm_a9_hps_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY        => arm_a9_hps_h2f_lw_axi_master_rready,  --                  .rready
			f2h_irq_p0           => arm_a9_hps_f2h_irq0_irq,              --          f2h_irq0.irq
			f2h_irq_p1           => arm_a9_hps_f2h_irq1_irq               --          f2h_irq1.irq
		);

	jtag_uart : component lab1_system_JTAG_UART
		port map (
			clk            => system_pll_sys_clk_clk,                                        --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	pushbuttons : component lab1_system_Pushbuttons
		port map (
			clk        => system_pll_sys_clk_clk,                           --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_1_pushbuttons_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_pushbuttons_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_pushbuttons_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_pushbuttons_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_pushbuttons_s1_readdata,        --                    .readdata
			in_port    => pushbuttons_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                          --                 irq.irq
		);

	system_pll : component lab1_system_System_PLL
		port map (
			ref_clk_clk        => system_pll_ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => system_pll_ref_reset_reset,    --    ref_reset.reset
			sys_clk_clk        => system_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => open,                          --    sdram_clk.clk
			reset_source_reset => system_pll_reset_source_reset  -- reset_source.reset
		);

	axi4_lite_count28_0 : component axi4_lite_count28
		generic map (
			C_S_AXI_DATA_WIDTH => 32,
			C_S_AXI_ADDR_WIDTH => 4
		)
		port map (
			clk                => system_pll_sys_clk_clk,                                  --     clock.clk
			reset_n            => rst_controller_reset_out_reset_ports_inv,                --     reset.reset_n
			out_leds           => leds_readdata,                                           --  out_leds.readdata
			axs_s0_AXI_AWADDR  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awaddr,  -- axi4_lite.awaddr
			axs_s0_AXI_AWPROT  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awprot,  --          .awprot
			axs_s0_AXI_AWVALID => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awvalid, --          .awvalid
			axs_s0_AXI_AWREADY => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awready, --          .awready
			axs_s0_AXI_WDATA   => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wdata,   --          .wdata
			axs_s0_AXI_WSTRB   => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wstrb,   --          .wstrb
			axs_s0_AXI_WVALID  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wvalid,  --          .wvalid
			axs_s0_AXI_WREADY  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wready,  --          .wready
			axs_s0_AXI_BRESP   => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bresp,   --          .bresp
			axs_s0_AXI_BVALID  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bvalid,  --          .bvalid
			axs_s0_AXI_BREADY  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bready,  --          .bready
			axs_s0_AXI_ARADDR  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_araddr,  --          .araddr
			axs_s0_AXI_ARPROT  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arprot,  --          .arprot
			axs_s0_AXI_ARVALID => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arvalid, --          .arvalid
			axs_s0_AXI_ARREADY => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arready, --          .arready
			axs_s0_AXI_RDATA   => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rdata,   --          .rdata
			axs_s0_AXI_RRESP   => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rresp,   --          .rresp
			axs_s0_AXI_RVALID  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rvalid,  --          .rvalid
			axs_s0_AXI_RREADY  => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rready   --          .rready
		);

	mm_interconnect_0 : component lab1_system_mm_interconnect_0
		port map (
			ARM_A9_HPS_h2f_axi_master_awid                                        => arm_a9_hps_h2f_axi_master_awid,                            --                                       ARM_A9_HPS_h2f_axi_master.awid
			ARM_A9_HPS_h2f_axi_master_awaddr                                      => arm_a9_hps_h2f_axi_master_awaddr,                          --                                                                .awaddr
			ARM_A9_HPS_h2f_axi_master_awlen                                       => arm_a9_hps_h2f_axi_master_awlen,                           --                                                                .awlen
			ARM_A9_HPS_h2f_axi_master_awsize                                      => arm_a9_hps_h2f_axi_master_awsize,                          --                                                                .awsize
			ARM_A9_HPS_h2f_axi_master_awburst                                     => arm_a9_hps_h2f_axi_master_awburst,                         --                                                                .awburst
			ARM_A9_HPS_h2f_axi_master_awlock                                      => arm_a9_hps_h2f_axi_master_awlock,                          --                                                                .awlock
			ARM_A9_HPS_h2f_axi_master_awcache                                     => arm_a9_hps_h2f_axi_master_awcache,                         --                                                                .awcache
			ARM_A9_HPS_h2f_axi_master_awprot                                      => arm_a9_hps_h2f_axi_master_awprot,                          --                                                                .awprot
			ARM_A9_HPS_h2f_axi_master_awvalid                                     => arm_a9_hps_h2f_axi_master_awvalid,                         --                                                                .awvalid
			ARM_A9_HPS_h2f_axi_master_awready                                     => arm_a9_hps_h2f_axi_master_awready,                         --                                                                .awready
			ARM_A9_HPS_h2f_axi_master_wid                                         => arm_a9_hps_h2f_axi_master_wid,                             --                                                                .wid
			ARM_A9_HPS_h2f_axi_master_wdata                                       => arm_a9_hps_h2f_axi_master_wdata,                           --                                                                .wdata
			ARM_A9_HPS_h2f_axi_master_wstrb                                       => arm_a9_hps_h2f_axi_master_wstrb,                           --                                                                .wstrb
			ARM_A9_HPS_h2f_axi_master_wlast                                       => arm_a9_hps_h2f_axi_master_wlast,                           --                                                                .wlast
			ARM_A9_HPS_h2f_axi_master_wvalid                                      => arm_a9_hps_h2f_axi_master_wvalid,                          --                                                                .wvalid
			ARM_A9_HPS_h2f_axi_master_wready                                      => arm_a9_hps_h2f_axi_master_wready,                          --                                                                .wready
			ARM_A9_HPS_h2f_axi_master_bid                                         => arm_a9_hps_h2f_axi_master_bid,                             --                                                                .bid
			ARM_A9_HPS_h2f_axi_master_bresp                                       => arm_a9_hps_h2f_axi_master_bresp,                           --                                                                .bresp
			ARM_A9_HPS_h2f_axi_master_bvalid                                      => arm_a9_hps_h2f_axi_master_bvalid,                          --                                                                .bvalid
			ARM_A9_HPS_h2f_axi_master_bready                                      => arm_a9_hps_h2f_axi_master_bready,                          --                                                                .bready
			ARM_A9_HPS_h2f_axi_master_arid                                        => arm_a9_hps_h2f_axi_master_arid,                            --                                                                .arid
			ARM_A9_HPS_h2f_axi_master_araddr                                      => arm_a9_hps_h2f_axi_master_araddr,                          --                                                                .araddr
			ARM_A9_HPS_h2f_axi_master_arlen                                       => arm_a9_hps_h2f_axi_master_arlen,                           --                                                                .arlen
			ARM_A9_HPS_h2f_axi_master_arsize                                      => arm_a9_hps_h2f_axi_master_arsize,                          --                                                                .arsize
			ARM_A9_HPS_h2f_axi_master_arburst                                     => arm_a9_hps_h2f_axi_master_arburst,                         --                                                                .arburst
			ARM_A9_HPS_h2f_axi_master_arlock                                      => arm_a9_hps_h2f_axi_master_arlock,                          --                                                                .arlock
			ARM_A9_HPS_h2f_axi_master_arcache                                     => arm_a9_hps_h2f_axi_master_arcache,                         --                                                                .arcache
			ARM_A9_HPS_h2f_axi_master_arprot                                      => arm_a9_hps_h2f_axi_master_arprot,                          --                                                                .arprot
			ARM_A9_HPS_h2f_axi_master_arvalid                                     => arm_a9_hps_h2f_axi_master_arvalid,                         --                                                                .arvalid
			ARM_A9_HPS_h2f_axi_master_arready                                     => arm_a9_hps_h2f_axi_master_arready,                         --                                                                .arready
			ARM_A9_HPS_h2f_axi_master_rid                                         => arm_a9_hps_h2f_axi_master_rid,                             --                                                                .rid
			ARM_A9_HPS_h2f_axi_master_rdata                                       => arm_a9_hps_h2f_axi_master_rdata,                           --                                                                .rdata
			ARM_A9_HPS_h2f_axi_master_rresp                                       => arm_a9_hps_h2f_axi_master_rresp,                           --                                                                .rresp
			ARM_A9_HPS_h2f_axi_master_rlast                                       => arm_a9_hps_h2f_axi_master_rlast,                           --                                                                .rlast
			ARM_A9_HPS_h2f_axi_master_rvalid                                      => arm_a9_hps_h2f_axi_master_rvalid,                          --                                                                .rvalid
			ARM_A9_HPS_h2f_axi_master_rready                                      => arm_a9_hps_h2f_axi_master_rready,                          --                                                                .rready
			System_PLL_sys_clk_clk                                                => system_pll_sys_clk_clk,                                    --                                              System_PLL_sys_clk.clk
			ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                        -- ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			JTAG_UART_reset_reset_bridge_in_reset_reset                           => rst_controller_reset_out_reset,                            --                           JTAG_UART_reset_reset_bridge_in_reset.reset
			JTAG_UART_avalon_jtag_slave_address                                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --                                     JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write                                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                                                .write
			JTAG_UART_avalon_jtag_slave_read                                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                                                .read
			JTAG_UART_avalon_jtag_slave_readdata                                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                                                .readdata
			JTAG_UART_avalon_jtag_slave_writedata                                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                                                .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest                               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                                                .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect                                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect   --                                                                .chipselect
		);

	mm_interconnect_1 : component lab1_system_mm_interconnect_1
		port map (
			ARM_A9_HPS_h2f_lw_axi_master_awid                                        => arm_a9_hps_h2f_lw_axi_master_awid,                       --                                       ARM_A9_HPS_h2f_lw_axi_master.awid
			ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      => arm_a9_hps_h2f_lw_axi_master_awaddr,                     --                                                                   .awaddr
			ARM_A9_HPS_h2f_lw_axi_master_awlen                                       => arm_a9_hps_h2f_lw_axi_master_awlen,                      --                                                                   .awlen
			ARM_A9_HPS_h2f_lw_axi_master_awsize                                      => arm_a9_hps_h2f_lw_axi_master_awsize,                     --                                                                   .awsize
			ARM_A9_HPS_h2f_lw_axi_master_awburst                                     => arm_a9_hps_h2f_lw_axi_master_awburst,                    --                                                                   .awburst
			ARM_A9_HPS_h2f_lw_axi_master_awlock                                      => arm_a9_hps_h2f_lw_axi_master_awlock,                     --                                                                   .awlock
			ARM_A9_HPS_h2f_lw_axi_master_awcache                                     => arm_a9_hps_h2f_lw_axi_master_awcache,                    --                                                                   .awcache
			ARM_A9_HPS_h2f_lw_axi_master_awprot                                      => arm_a9_hps_h2f_lw_axi_master_awprot,                     --                                                                   .awprot
			ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     => arm_a9_hps_h2f_lw_axi_master_awvalid,                    --                                                                   .awvalid
			ARM_A9_HPS_h2f_lw_axi_master_awready                                     => arm_a9_hps_h2f_lw_axi_master_awready,                    --                                                                   .awready
			ARM_A9_HPS_h2f_lw_axi_master_wid                                         => arm_a9_hps_h2f_lw_axi_master_wid,                        --                                                                   .wid
			ARM_A9_HPS_h2f_lw_axi_master_wdata                                       => arm_a9_hps_h2f_lw_axi_master_wdata,                      --                                                                   .wdata
			ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       => arm_a9_hps_h2f_lw_axi_master_wstrb,                      --                                                                   .wstrb
			ARM_A9_HPS_h2f_lw_axi_master_wlast                                       => arm_a9_hps_h2f_lw_axi_master_wlast,                      --                                                                   .wlast
			ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      => arm_a9_hps_h2f_lw_axi_master_wvalid,                     --                                                                   .wvalid
			ARM_A9_HPS_h2f_lw_axi_master_wready                                      => arm_a9_hps_h2f_lw_axi_master_wready,                     --                                                                   .wready
			ARM_A9_HPS_h2f_lw_axi_master_bid                                         => arm_a9_hps_h2f_lw_axi_master_bid,                        --                                                                   .bid
			ARM_A9_HPS_h2f_lw_axi_master_bresp                                       => arm_a9_hps_h2f_lw_axi_master_bresp,                      --                                                                   .bresp
			ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      => arm_a9_hps_h2f_lw_axi_master_bvalid,                     --                                                                   .bvalid
			ARM_A9_HPS_h2f_lw_axi_master_bready                                      => arm_a9_hps_h2f_lw_axi_master_bready,                     --                                                                   .bready
			ARM_A9_HPS_h2f_lw_axi_master_arid                                        => arm_a9_hps_h2f_lw_axi_master_arid,                       --                                                                   .arid
			ARM_A9_HPS_h2f_lw_axi_master_araddr                                      => arm_a9_hps_h2f_lw_axi_master_araddr,                     --                                                                   .araddr
			ARM_A9_HPS_h2f_lw_axi_master_arlen                                       => arm_a9_hps_h2f_lw_axi_master_arlen,                      --                                                                   .arlen
			ARM_A9_HPS_h2f_lw_axi_master_arsize                                      => arm_a9_hps_h2f_lw_axi_master_arsize,                     --                                                                   .arsize
			ARM_A9_HPS_h2f_lw_axi_master_arburst                                     => arm_a9_hps_h2f_lw_axi_master_arburst,                    --                                                                   .arburst
			ARM_A9_HPS_h2f_lw_axi_master_arlock                                      => arm_a9_hps_h2f_lw_axi_master_arlock,                     --                                                                   .arlock
			ARM_A9_HPS_h2f_lw_axi_master_arcache                                     => arm_a9_hps_h2f_lw_axi_master_arcache,                    --                                                                   .arcache
			ARM_A9_HPS_h2f_lw_axi_master_arprot                                      => arm_a9_hps_h2f_lw_axi_master_arprot,                     --                                                                   .arprot
			ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     => arm_a9_hps_h2f_lw_axi_master_arvalid,                    --                                                                   .arvalid
			ARM_A9_HPS_h2f_lw_axi_master_arready                                     => arm_a9_hps_h2f_lw_axi_master_arready,                    --                                                                   .arready
			ARM_A9_HPS_h2f_lw_axi_master_rid                                         => arm_a9_hps_h2f_lw_axi_master_rid,                        --                                                                   .rid
			ARM_A9_HPS_h2f_lw_axi_master_rdata                                       => arm_a9_hps_h2f_lw_axi_master_rdata,                      --                                                                   .rdata
			ARM_A9_HPS_h2f_lw_axi_master_rresp                                       => arm_a9_hps_h2f_lw_axi_master_rresp,                      --                                                                   .rresp
			ARM_A9_HPS_h2f_lw_axi_master_rlast                                       => arm_a9_hps_h2f_lw_axi_master_rlast,                      --                                                                   .rlast
			ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      => arm_a9_hps_h2f_lw_axi_master_rvalid,                     --                                                                   .rvalid
			ARM_A9_HPS_h2f_lw_axi_master_rready                                      => arm_a9_hps_h2f_lw_axi_master_rready,                     --                                                                   .rready
			axi4_lite_count28_0_axi4_lite_awaddr                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awaddr,  --                                      axi4_lite_count28_0_axi4_lite.awaddr
			axi4_lite_count28_0_axi4_lite_awprot                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awprot,  --                                                                   .awprot
			axi4_lite_count28_0_axi4_lite_awvalid                                    => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awvalid, --                                                                   .awvalid
			axi4_lite_count28_0_axi4_lite_awready                                    => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_awready, --                                                                   .awready
			axi4_lite_count28_0_axi4_lite_wdata                                      => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wdata,   --                                                                   .wdata
			axi4_lite_count28_0_axi4_lite_wstrb                                      => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wstrb,   --                                                                   .wstrb
			axi4_lite_count28_0_axi4_lite_wvalid                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wvalid,  --                                                                   .wvalid
			axi4_lite_count28_0_axi4_lite_wready                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_wready,  --                                                                   .wready
			axi4_lite_count28_0_axi4_lite_bresp                                      => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bresp,   --                                                                   .bresp
			axi4_lite_count28_0_axi4_lite_bvalid                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bvalid,  --                                                                   .bvalid
			axi4_lite_count28_0_axi4_lite_bready                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_bready,  --                                                                   .bready
			axi4_lite_count28_0_axi4_lite_araddr                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_araddr,  --                                                                   .araddr
			axi4_lite_count28_0_axi4_lite_arprot                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arprot,  --                                                                   .arprot
			axi4_lite_count28_0_axi4_lite_arvalid                                    => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arvalid, --                                                                   .arvalid
			axi4_lite_count28_0_axi4_lite_arready                                    => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_arready, --                                                                   .arready
			axi4_lite_count28_0_axi4_lite_rdata                                      => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rdata,   --                                                                   .rdata
			axi4_lite_count28_0_axi4_lite_rresp                                      => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rresp,   --                                                                   .rresp
			axi4_lite_count28_0_axi4_lite_rvalid                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rvalid,  --                                                                   .rvalid
			axi4_lite_count28_0_axi4_lite_rready                                     => mm_interconnect_1_axi4_lite_count28_0_axi4_lite_rready,  --                                                                   .rready
			System_PLL_sys_clk_clk                                                   => system_pll_sys_clk_clk,                                  --                                                 System_PLL_sys_clk.clk
			ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                      -- ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			axi4_lite_count28_0_reset_reset_bridge_in_reset_reset                    => rst_controller_reset_out_reset,                          --                    axi4_lite_count28_0_reset_reset_bridge_in_reset.reset
			Pushbuttons_reset_reset_bridge_in_reset_reset                            => rst_controller_001_reset_out_reset,                      --                            Pushbuttons_reset_reset_bridge_in_reset.reset
			Pushbuttons_s1_address                                                   => mm_interconnect_1_pushbuttons_s1_address,                --                                                     Pushbuttons_s1.address
			Pushbuttons_s1_write                                                     => mm_interconnect_1_pushbuttons_s1_write,                  --                                                                   .write
			Pushbuttons_s1_readdata                                                  => mm_interconnect_1_pushbuttons_s1_readdata,               --                                                                   .readdata
			Pushbuttons_s1_writedata                                                 => mm_interconnect_1_pushbuttons_s1_writedata,              --                                                                   .writedata
			Pushbuttons_s1_chipselect                                                => mm_interconnect_1_pushbuttons_s1_chipselect              --                                                                   .chipselect
		);

	irq_mapper : component lab1_system_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq, -- receiver1.irq
			sender_irq    => arm_a9_hps_f2h_irq0_irq   --    sender.irq
		);

	irq_mapper_001 : component lab1_system_irq_mapper_001
		port map (
			clk        => open,                    --       clk.clk
			reset      => open,                    -- clk_reset.reset
			sender_irq => arm_a9_hps_f2h_irq1_irq  --    sender.irq
		);

	rst_controller : component lab1_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,        -- reset_in1.reset
			clk            => system_pll_sys_clk_clk,               --       clk.clk
			reset_out      => rst_controller_reset_out_reset,       -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_001 : component lab1_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => system_pll_reset_source_reset,      -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component lab1_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,               --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_in1      => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_1_pushbuttons_s1_write_ports_inv <= not mm_interconnect_1_pushbuttons_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	arm_a9_hps_h2f_reset_reset_ports_inv <= not arm_a9_hps_h2f_reset_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of lab1_system
