
module lab (
	);	

endmodule
